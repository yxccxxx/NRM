IEEE round to nearest, even on tie

1.4999999999 ==> 1
1.5 ==> 2
1.50000000001 ==> 2

2.4999999999 ==> 2
2.5 ==> 2
2.50000000001 ==> 3

1??_????_????_????	  2**14

1.???????????  2**0

exp = 29 = 14 + bias = 14 + 15

111_1111_1111_1111  2**15-1
1.111111111111 1.11111 * 2**14